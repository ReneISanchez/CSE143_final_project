------------------------------------------------------------------------------
-- i2c slave receiver
------------------------------------------------------------------------------
-- Intended target: Xilinx CoolRunner-II CPLD  (XC2C64A)
-- Development tools: XILINX ISE 7.1i webpack
-- Author:  DMITRY PETROV
-- Notes:
-- Date:     11-09-2005
-- Revision: 1.0
------------------------------------------------------------------------------
-- This code implements i2c slave which is able to receive a data byte.
 
-- i2c message has 3 parts:
-- <Device Address> 22h
-- <Sub Address> 00h
-- <Data byte> XX 
-- If Device and Sub Addresses are matched the data byte will be accepted.

-- Because of SCL line used as clock for i2c state machine, slow SCL changes 
-- will make noise and invalid data reception. 

-- To avoid noise of slow SCL - usualy used an external CLOCK, for 
-- clocking all modules but it will take some amount of CPLD's macrocells.

-- Another way is to use an SCHMITT TRIGGER on SCL and SDA. 
-- Forexample XILINX CoolRunner-II CPLD, has SCHMITT TRIGGER on it's I/O.
-- By default this function is deactivated, PLEASE ACTIVATE IT !

-- If your PLD have no SCHMITT TRIGGER function, you may use solution wich 
-- require 2 resistors and aditional output pin. 
-- Here's an old Xilinx app note about it: 
-- http://www.xilinx.com/xcell/xl19/xl19-34.pdf 
-- ===========================================================================
-- DISCLAIMER: This code is FREEWARE which is provided on an �as is� basis, 
-- YOU MAY USE IT ON YOUR OWN RISK, WITHOUT ANY WARRANTY. 
-- ===========================================================================d

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

------------------------------------------------------------------------------
entity i2c_m_rx is
	generic(
		DADDR		: std_logic_vector(6 downto 0) := "0000001";		   -- 11h (22h) device address
		ADDR		: std_logic_vector(7 downto 0)  := "00000000"		   -- 00h	    sub address		
	);
	port(
		CLK		: in std_logic;
		RST		: in std_logic;
		SCL		: out std_logic := '0';
		SDA		: inout std_logic;
		DIN 		: in std_logic_vector(7 downto 0);			   -- Recepted over i2c data byte
		DOUT 		: out std_logic_vector(7 downto 0) := "00000000"
	);
	--SCHMITT TRIGGER activation (folowing 3 strings should be uncommented)
	--attribute SCHMITT_TRIGGER: string; 
	--attribute SCHMITT_TRIGGER of SCL: signal is "true"; 
	--attribute SCHMITT_TRIGGER of SDA: signal is "true";
end i2c_m_rx;

------------------------------------------------------------------------------
architecture Behavioral of i2c_m_rx is
	signal DOUT_S: std_logic_vector(7 downto 0);
	signal SDA_IN, START, START_RST, STOP, ACTIVE, ACK	: std_logic;
	signal SHIFTREG	: std_logic_vector(8 downto 0) := "000000000";
	signal STATE : std_logic_vector(1 downto 0) := "00";		-- 00 - iddle state	
	signal addrData : std_logic;																		-- 01 - DADDR  compare
	signal count : std_logic_vector(3 downto 0);
	signal reset : std_logic;-- 10 - ADDR compare	-- 11 - DATA read
	signal scl_val : std_logic := '0';
begin

process (CLK)
begin 
	if(CLK'EVENT and CLK = '1') then
			SCL <= '1';
			scl_val <= '1';
	elsif(CLK'EVENT and CLK = '0') then  
			SCL <= '0';
			scl_val <= '0';
	end if;
end process;

-- stop condition detection
process (RST, scl_val, SDA, START, reset)
begin
	if (RST = '0' or (scl_val = '0')) or START = '1' or reset = '0' then
		STOP <= '0';
		reset <= '1';
		if(STATE = "00") then
			addrData <= '0';
			count <= "0110";
		end if;
	elsif scl_val = '1' and (SDA = '1' and SDA'EVENT) then
		STOP <= '1';
	end if;
end process;

------------------------------------------------------------------------------
-- start condition detection, method 2 ( simple - but week against noise )
process (RST, scl_val, SDA_IN, START)
begin
	if (SDA = '0' and (scl_val = '0' and scl_val'EVENT))  then
		START <= '1';
		if(STATE = "01") then
			count <= "0111";
		end if;
	elsif scl_val = '1' and (SDA = '0' and SDA'event) then
		START <= '0';
	end if;
end process;

------------------------------------------------------------------------------
-- "active communication" signal 
process (RST, STOP, START)
begin
	if RST = '0' or STOP = '1' then	 --or (SHIFTREG="000000001" and ACK = '0' and SCL='1' and SCL'event) 
		ACTIVE <= '0';
	elsif START = '0' and START'event then
		ACTIVE <= '1';
	end if;
end process;

------------------------------------------------------------------------------
-- WX data shifter
process (RST, ACTIVE, ACK, scl_val, SDA_IN)
begin 
if (STATE = "10" or STATE = "01") and (scl_val = '1' and scl_val'EVENT) then
	if(SDA = '0') then
		DOUT <= "11111111";
		addrData <= '1';
		STATE <= "11";
	else 
		DOUT <= "00000000";
	end if;
	--SHIFTREG <= "000000001";	

		--SHIFTREG(8 downto 0) <= SHIFTREG(7 downto 0) & SDA_IN;
end if;							  
end process;

------------------------------------------------------------------------------
-- I2C data write
process (RST, SHIFTREG, addrData, START, STATE,count)
begin
if RST = '0' then
	DOUT_S <= "00000000";
elsif addrData='0' and (START = '0' and START'EVENT) and (count /= "1111") then	
	SDA <= DADDR(to_integer(unsigned (count)));
	count <= std_logic_vector(unsigned(count) - "0001");
	STATE <= "00";
elsif count = "1111" and addrData = '0'  then
	SDA <= '0';
	STATE <= "01";
elsif count >= "0000" and addrData = '1' and (START = '0' and START'EVENT) then
	SDA <= DIN(to_integer(unsigned(count)));
	count <= std_logic_vector(unsigned(count) - "0001");
   if count = "0000" then
		STATE <= "10";
	end if;
elsif addrData = '1' and STATE = "11" then
	reset <= '0';
	STATE <= "00";
	addrData <= '0';
end if;
end process; 

------------------------------------------------------------------------------
--DIN(7 downto 0) <= DOUT_S(7 downto 0);

end Behavioral;
------------------------------------------------------------------------------